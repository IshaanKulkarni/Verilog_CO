module addsub(a,b,c,d,e);
input reg [31:0]a;
input reg [31:0]b;
input c;
output [31:0]d;
output [31:0]e;
wire [31:0]s;
if(c==1)



end

endmodule