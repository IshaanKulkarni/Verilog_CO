module func_testbench;
reg [31:0]A;
reg [31:0]B;
reg [31:0]C;
reg [31:0]D;
reg [31:0]E;
reg [31:0]F;
wire[31:0]AN;
wire[31:0]OR;
wire[31:0]NOR;
and18 Ishaandut18(.c(AN),.a(A),.b(B));
or18 Ishaandut19(.f(OR),.d(C),.e(D));
nor18 Ishaandut20(.j(NOR),.g(E),.h(F));
initial
begin
A = 'b00100100001100110011001010101010; B = 'b10101100110010101010101010101010; C='b10101111111111110000110011001100; D='b10101111111111111111111111111111; E='b01010000000000000000000000000101; F='b00101011111111110000000010101010 ;
#10 A ='b01011110101000000011000010101010; B = 'b11111111111111110010101010101010; C='b10101010101010101010101010101010; D='b10101111110101010101010101010111; E='b10101010111111111111111111110101; F='b10111010101010101010111111000011;

end

endmodule