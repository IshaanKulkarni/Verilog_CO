module ALUTB;
reg [31:0]A;
reg [31:0]B;
reg [32:0]C;
reg s0,s1,s2;

ALU dut_Ishaan(.res(C),.a(A),.b(B),.s0(s0),.s1(s1),.s2(s2));
initial
begin
A = 'b10101010100001010101010; B = 'b0111011101010010; s2=0;s1=0;s0=0;  
#100 A = 'b10101010101010101010101010001000; B = 'b10100010100010; s2=0;s1=0;s0=0;
#100 A = 'b10100010001010000000010010101011; B = 'b00100101010010; s2=0;s1=1;s0=0;
#100 A = 'b10001010000010001010000010101100; B = 'b10100010001010; s2=0;s1=1;s0=1;
end

endmodule