module rca_testbench;
reg [31:0]A;
reg [31:0]B;
reg Cin;
wire [31:0]S,C;
rca Ishaan_dut(.sum(S),.cout(C),.a(A),.b(B),.cin(Cin));
initial
begin
A = 'b00000000000000000000000000000000; B = 'b001111111111111111111111111111; Cin=0; 
#10 A = 'b01010101010101010101010101010101; B = 'b111111111111111111111111111111; Cin=0;
#10 A = 'b10101010101010101011100010101101; B = 'b011011011011100011101010011001; Cin=0;
#10 A = 'b11111111111111111111111111111001; B = 'b101000001000100001010000100010; Cin=0;
end

endmodule